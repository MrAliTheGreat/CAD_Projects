library verilog;
use verilog.vl_types.all;
entity TestBenchRecursive is
end TestBenchRecursive;
