library verilog;
use verilog.vl_types.all;
entity INV_gate is
    port(
        \out\           : out    vl_logic;
        in1             : in     vl_logic
    );
end INV_gate;
