library verilog;
use verilog.vl_types.all;
entity TB_Circuit is
end TB_Circuit;
