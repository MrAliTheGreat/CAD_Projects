library verilog;
use verilog.vl_types.all;
entity StackTestBench is
end StackTestBench;
