library verilog;
use verilog.vl_types.all;
entity MemoriesTestBench is
end MemoriesTestBench;
